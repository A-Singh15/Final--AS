module accumulator (
    output  reg  [15:0] sum,  // accumulated out
    input   [7:0]       in,   // input
    input               rst,  // reset
    input               clk   // clock
);
    wire carry;
    wire [15:0] sum_in;
    
    assign {carry, sum_in} = sum + in;
    
    always @(posedge clk) begin
        if (rst) begin
            sum <= 0;
        end else begin
            sum <= (carry) ? 16'hFFFF : sum_in;
        end
    end
endmodule
